LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.PIPELINE.ALL;
USE WORK.TOOLBOX.ALL;

ENTITY DUMMY IS 
	
	GENERIC ( CTRL_WORD_TOTAL : INTEGER := 20; CTRL_WORD_OUT : INTEGER := 18);
	PORT 	( 	
				CLK,RST    : IN  STD_LOGIC;						--\
				WB_RD_LOAD : IN  STD_LOGIC_VECTOR(4  DOWNTO 0); --| Register File inputs.
				WB_RD_DATA : IN  STD_LOGIC_VECTOR(31 DOWNTO 0); --/ 	
				PC_VALUE   : IN  STD_LOGIC_VECTOR(31 DOWNTO 0); -- Feed from
				IF_WORD    : IN  STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction Fetch
				
				RD_FROM_EXE: IN  STD_LOGIC_VECTOR(4  DOWNTO 0);
				RD_FROM_MEM: IN  STD_LOGIC_VECTOR(4  DOWNTO 0);
				PIPE_LOAD_E: IN  STD_LOGIC;

				RS1_VALUE  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); 
				RS2_VALUE  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				RD_ADDR    : OUT STD_LOGIC_VECTOR(4  DOWNTO 0);
				IMMEDIATE  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				TARGET_AD  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); 
				PC_VALUE_O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				CTRL_WORD  : OUT STD_LOGIC_VECTOR(CTRL_WORD_OUT-1  DOWNTO 0);
				
				PIPE_STALL : OUT STD_LOGIC;
				PIPE_FWDA  : OUT STD_LOGIC_VECTOR(1 DOWNTO 0); 
				PIPE_FWDB  : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
				PIPE_FWDC  : OUT STD_LOGIC

			);

END DUMMY;


ARCHITECTURE ULTRA_DUMMY OF DUMMY IS;
	
	
	BEGIN
	
	ID2: I_D
		 GENERIC MAP( CTRL_WORD_TOTAL => 20, CTRL_WORD_OUT => 18 )
		 PORT    MAP(	
						CLK 	   => CLK,
						RST 	   => RST,
						WB_RD_LOAD => ID_IN_WB_RD_ADR, -- Input from WB
						WB_RD_DATA => ID_IN_WB_RD_VAL, -- Input from S
						PC_VALUE   => PIPE_OUT_PC_VAL, -- 
						IF_WORD    => PIPE_OUT_IFWORD, -- 
						RD_FROM_EXE=> ID_IN_RD_EXE,
						RD_FROM_MEM=> ID_IN_RD_MEM,
						PIPE_LOAD_E=> ID_IN_LOAD_EXE,
						RS1_VALUE  => ID_OUT_RS1_VAL,
						RS2_VALUE  => ID_OUT_RS2_VAL,
						RD_ADDR    => ID_OUT_RD_ADR,
						IMMEDIATE  => ID_OUT_IMM,
						TARGED_AD  => ID_OUT_J_TARGET,
						PC_VALUE_O => ID_OUT_PC_VAL,
						CTRL_WORD  => ID_OUT_OPCODES,
						PIPE_STALL => PIPE_STALL_SIG,
						PIPE_FWDA  => ID_OUT_FWD_A,
						PIPE_FWDB  => ID_OUT_FWD_B,
						PIPE_FWDC  => ID_OUT_FWDC
					);
END ULTRA_DUMMY;
