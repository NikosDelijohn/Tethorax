-- Casual 32 to 1 Generic input Multiplexer.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX32X1 IS

	GENERIC( INSIZE : INTEGER := 10 );
	
	PORT(
	
			D0 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D1 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D2 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D3 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D4 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D5 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D6 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D7 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D8 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D9 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D10: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D11: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D12: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D13: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D14: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D15: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D16: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D17: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D18: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D19: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D20: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D21: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D22: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D23: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D24: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D25: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D26: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D27: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D28: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D29: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D30: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D31: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			
			SEL: IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
			
			O  : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
	    );
		
END MUX32X1;

ARCHITECTURE RTL OF MUX32X1 IS

BEGIN

	PROCESS(SEL,D0 ,D1 ,D2 ,D3 ,D4 ,D5 ,D6 ,D7 ,D8 ,D9 ,D10,D11,D12,D13,D14,D15,
	            D16,D17,D18,D19,D20,D21,D22,D23,D24,D25,D26,D27,D28,D29,D30,D31)
	BEGIN
	
		CASE SEL IS
		    	--    OPCODE
			WHEN "00000" => O <= D0;  -- LOADS
			WHEN "00001" => O <= D1;  
			WHEN "00010" => O <= D2;
			WHEN "00011" => O <= D3;
			WHEN "00100" => O <= D4;  -- I-OPS
			WHEN "00101" => O <= D5;  -- AUIPC
			WHEN "00110" => O <= D6;
			WHEN "00111" => O <= D7;
			WHEN "01000" => O <= D8;  -- STORES
			WHEN "01001" => O <= D9;
			WHEN "01010" => O <= D10;
			WHEN "01011" => O <= D11;
			WHEN "01100" => O <= D12; -- R-OPS
			WHEN "01101" => O <= D13; -- LUI
			WHEN "01110" => O <= D14;
			WHEN "01111" => O <= D15;
			WHEN "10000" => O <= D16;
			WHEN "10001" => O <= D17;
			WHEN "10010" => O <= D18;
			WHEN "10011" => O <= D19;
			WHEN "10100" => O <= D20;
			WHEN "10101" => O <= D21;
			WHEN "10110" => O <= D22;
			WHEN "10111" => O <= D23;
			WHEN "11000" => O <= D24; -- BRANCHES
			WHEN "11001" => O <= D25; -- JALR
			WHEN "11010" => O <= D26;
			WHEN "11011" => O <= D27; -- JAL
			WHEN "11100" => O <= D28;
			WHEN "11101" => O <= D29;
			WHEN "11110" => O <= D30;
			WHEN "11111" => O <= D31;
			WHEN OTHERS  => O <= (OTHERS => 'X');
		
		END CASE;
		
	END PROCESS;
	
END RTL;
