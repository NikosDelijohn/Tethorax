LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY PC_PLUS_4 IS

	PORT (
			PC : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
			RES: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		 );

END PC_PLUS_4;

ARCHITECTURE BEHAVIORAL OF PC_PLUS_4 IS
	
	SIGNAL FOUR : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000100";
	BEGIN
	
	RES <= STD_LOGIC_VECTOR(UNSIGNED(PC) + UNSIGNED(FOUR));
	
END BEHAVIORAL;