-- This is a Custom PACKAGE file used to avoid duplicate code being written
-- in other files (e.g. ARCHITECTURES).

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE TOOLBOX IS

-- ================== INSTRUCTION FETCH COMPONENTS ================== --
------------------------------------------------------------------------
	-- Defined @ "I_F_RAM.vhd" file.
	COMPONENT I_F_RAM IS
	
			PORT
				(
					address		: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
					clock		: IN STD_LOGIC  := '1';
					data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
					wren		: IN STD_LOGIC ;
					q		    : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
				);
				
	END COMPONENT I_F_RAM;
	
-- ================== INSTRUCTION DECODE COMPONENTS ================== --
-------------------------------------------------------------------------
	-- Defined @ "MUX2X1.vhd" file.
	COMPONENT MUX2X1 IS

		GENERIC ( INSIZE : INTEGER := 10 );
	
		PORT (
				A : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				B : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			  SEL : IN  STD_LOGIC;
				O : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
			 );

	END COMPONENT MUX2X1;
	
-------------------------------------------------------------------------
	-- Defined @ "MUX8X1.vhd" file.
	COMPONENT MUX8X1 IS 
		-- Defined @ "MUX8X1.vhd" file.
		GENERIC ( INSIZE : INTEGER := 10 );
		
		PORT (	
				D0  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D1  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D2  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D3  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D4  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D5  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D6  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D7  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				
				SEL : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
			 
				O : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
			 );

	END COMPONENT MUX8X1;
-------------------------------------------------------------------------
	-- Defined @ "MUX32X1.vhd" file.
	COMPONENT MUX32X1 IS

		GENERIC ( INSIZE : INTEGER := 10 );
		
		PORT (
		
				 D0: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D1: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D2: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D3: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D4: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D5: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D6: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D7: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D8: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				 D9: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D10: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D11: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D12: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D13: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D14: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D15: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D16: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D17: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D18: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D19: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D20: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D21: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D22: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D23: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D24: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D25: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D26: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D27: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D28: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D29: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D30: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				D31: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
				
				SEL: IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
				
				O  : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
			);
			
	END COMPONENT MUX32X1;
-------------------------------------------------------------------------	
END PACKAGE TOOLBOX;