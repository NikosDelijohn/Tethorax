
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


USE WORK.PIPELINE.ALL;
USE WORK.TOOLBOX.ALL;

ENTITY ASDF IS
	PORT( A: IN BIT;
          B: OUT BIT);
END ASDF;

ARCHITECTURE E OF ASDF IS

	SIGNAL ID_IN_WB_RD_ADR: STD_LOGIC_VECTOR(4  DOWNTO 0);
	SIGNAL ID_IN_WB_RD_VAL: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_IN_RD_EXE   : STD_LOGIC_VECTOR(4  DOWNTO 0);
	SIGNAL ID_IN_RD_MEM   : STD_LOGIC_VECTOR(4  DOWNTO 0);
	SIGNAL ID_IN_LOAD_EXE : STD_LOGIC;
	SIGNAL ID_OUT_RS1_VAL : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_OUT_RS2_VAL : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_OUT_RD_ADR  : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL ID_OUT_IMM     : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_OUT_J_TARGET: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_OUT_PC_VAL  : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_OUT_OPCODES : STD_LOGIC_VECTOR(17 DOWNTO 0);
	SIGNAL ID_OUT_STALL   : STD_LOGIC;
	SIGNAL ID_OUT_FWD_A   : STD_LOGIC_VECTOR(1  DOWNTO 0);
	SIGNAL ID_OUT_FWD_B   : STD_LOGIC_VECTOR(1  DOWNTO 0);
	SIGNAL ID_OUT_FWD_C   : STD_LOGIC;
	SIGNAL PIPE_STALL_SIG : STD_LOGIC;
	
	SIGNAL CLK: STD_LOGIC;
	SIGNAL RST:STD_LOGIC;
	
	signal ID_OUT_RS1_VALe : std_logic_vector(31 downto 0);
	signal ID_OUT_RS1_VALb : std_logic_vector(31 downto 0);
	
	BEGIN 

	ID2: I_D
		 GENERIC MAP( CTRL_WORD_TOTAL => 20, CTRL_WORD_OUT => 18 )
		 PORT    MAP(	
						CLK 	   => CLK,
						RST 	   => RST,
						WB_RD_LOAD => ID_IN_WB_RD_ADR, -- Input from WB
						WB_RD_DATA => ID_IN_WB_RD_VAL, -- Input from S
						PC_VALUE   => ID_OUT_RS1_VALe, -- 
						IF_WORD    => ID_OUT_RS1_VALb, -- 
						RD_FROM_EXE=> ID_IN_RD_EXE,
						RD_FROM_MEM=> ID_IN_RD_MEM,
						PIPE_LOAD_E=> ID_IN_LOAD_EXE,
						RS1_VALUE  => ID_OUT_RS1_VAL,
						RS2_VALUE  => ID_OUT_RS2_VAL,
						RD_ADDR    => ID_OUT_RD_ADR,
						IMMEDIATE  => ID_OUT_IMM,
						TARGET_AD  => ID_OUT_J_TARGET,
						PC_VALUE_O => ID_OUT_PC_VAL,
						CTRL_WORD  => ID_OUT_OPCODES,
						PIPE_STALL => PIPE_STALL_SIG,
						PIPE_FWDA  => ID_OUT_FWD_A,
						PIPE_FWDB  => ID_OUT_FWD_B,
						PIPE_FWDC  => ID_OUT_FWD_C
					);

END E;