-- Casual 2x1 Mux of STD_LOGIC type

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX2X1_BIT IS

	PORT ( 
			D0  : IN  STD_LOGIC;
			D1  : IN  STD_LOGIC;
		    SEL : IN  STD_LOGIC;
		    O   : OUT STD_LOGIC
		 );
		 
END MUX2X1_BIT;

ARCHITECTURE BEHAVIORAL OF MUX2X1_BIT IS

	BEGIN
	
	O <= D0 WHEN (SEL = '0') ELSE D1;
	
END BEHAVIORAL;