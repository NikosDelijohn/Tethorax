-- Structural Component on which the 32bit Adder/Subber is based on

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXE_ADDER_SUBBER_CELL IS 

	PORT(
		A  : IN  STD_LOGIC; 
		B  : IN  STD_LOGIC;
		CI : IN  STD_LOGIC;
		OP : IN  STD_LOGIC; -- O = ADD / 1 = INVERT B
		S  : OUT STD_LOGIC;
		CO : OUT STD_LOGIC
	    );
		 
END EXE_ADDER_SUBBER_CELL;

ARCHITECTURE RTL OF EXE_ADDER_SUBBER_CELL IS 

	SIGNAL B_XOR_MODE  : STD_LOGIC;
	SIGNAL PARTIAL_SUM : STD_LOGIC;
	
	BEGIN 
	
	B_XOR_MODE  <= B XOR OP;
	
	PARTIAL_SUM <= B_XOR_MODE XOR A;
	CO          <= (A AND B_XOR_MODE) OR ( PARTIAL_SUM AND CI);
	S 	    <= PARTIAL_SUM XOR CI;
	
	
END RTL;