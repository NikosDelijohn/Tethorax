-- Typical 8 to 1 Generic input Multiplexer.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX8X1 IS 
	
	GENERIC ( INSIZE : INTEGER := 10 );
	
	PORT (	
			D0  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D1  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D2  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D3  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D4  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D5  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D6  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D7  : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			
		    SEL : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		 
		    O : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
		 );

END MUX8X1;

ARCHITECTURE RTL OF MUX8X1 IS
BEGIN
	PROCESS(SEL)
	BEGIN
		CASE SEL IS 
		
			WHEN "000" => O <= D0;
			WHEN "001" => O <= D1;
			WHEN "010" => O <= D2;
			WHEN "011" => O <= D3;
			WHEN "100" => O <= D4;
			WHEN "101" => O <= D5;
			WHEN "110" => O <= D6;
			WHEN "111" => O <= D7;
			
			WHEN OTHERS => O <= (OTHERS =>'Z');
			
		END CASE;
	END PROCESS;
	
END RTL;