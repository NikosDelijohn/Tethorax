LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REG_FLIPPER IS

	PORT (
			IF_WORD : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
			FLIP    : OUT STD_LOGIC
		 );
		 
END REG_FLIPPER;

ARCHITECTURE RTL OF REG_FLIPPER IS

	SIGNAL BGE  : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL BGEU : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RES  : STD_LOGIC_VECTOR(2 DOWNTO 0);
		
	BEGIN
	
	BGE  <= "101";
	BGEU <= "111";
	
	RES  <= ( BGE XNOR IF_WORD) OR ( BGEU XNOR IF_WORD);
	FLIP <= RES(0) AND RES(1) AND RES(2);
	
END RTL;
