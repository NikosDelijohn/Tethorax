LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDER_2B IS

	PORT ( 
			A  : IN STD_LOGIC;
			B  : IN STD_LOGIC;
			CI : IN STD_LOGIC;
			S  : OUT STD_LOGIC;
			CO : OUT STD_LOGIC 
		 );

END ADDER_2B;

ARCHITECTURE RTL OF ADDER_2B IS

	SIGNAL PARTIAL_SUM : STD_LOGIC;

	BEGIN 

		PARTIAL_SUM <= A XOR B;
		S			<= PARTIAL_SUM XOR CI;
		CO			<= (A AND B) OR (CI AND PARTIAL_SUM);

END RTL;