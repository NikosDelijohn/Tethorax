LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;

USE WORK.TOOLBOX.ALL;

ENTITY MEM_TO_WB IS

	PORT(
		  MEM_IN: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		  ALU_IN: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		  MEMOP : IN  STD_LOGIC_VECTOR(2  DOWNTO 0);

		  WB_IN : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	    );

END MEM_TO_WB;

ARCHITECTURE STRUCTURAL OF MEM_TO_WB IS

	SIGNAL MUX_SEL : STD_LOGIC;
	
	BEGIN

	MUX_SEL <= AND_REDUCE(MEMOP);

	MUX: MUX2X1
		 GENERIC MAP ( INSIZE => 32 )
		 PORT    MAP (
					   D0  => MEM_IN,
					   D1  => ALU_IN,
					   SEL => MUX_SEL,
					   O   => WB_IN
					 );

END STRUCTURAL;