
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY WORK;
USE WORK.TOOLBOX.ALL;

ENTITY REGISTER_FILE IS 

	PORT ( 
			CLK,RST  : IN STD_LOGIC;
			LOAD_REG : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		    ADDR_RS1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			ADDR_RS2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := NULL;
			DATA_IN  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		 );
		 
END REGISTER_FILE;

ARCHITECTURE STRUCTURAL OF REGISTER_FILE IS
	
	TYPE MATRIX_2D IS ARRAY (0 TO 31, 31 DOWNTO 0) OF STD_LOGIC_VECTOR;
	
	SIGNAL BUF_OF_BUFFERS : MATRIX_2D(0 TO 31, 31 DOWNTO 0);
	
	BEGIN 
	
		GEN: FOR I IN 0 TO 31 GENERATE 
		
			CASE0: IF I = 0 GENERATE
				   
				   ZERO_REG: REG_32B_ZERO
							 PORT MAP( 
									   CLK => CLK,
									   Q_OUT => BUF_OF_BUFFERS(I,31 DOWNTO 0) -- <== PROBLEM HERE.
							         );
			END GENERATE CASE0;
							         
			CASE1: IF I > 0 AND I <= 31 GENERATE
				   
				   CASUALS:  REG_32B_CASUAL
							 PORT MAP(
										LOAD  => LOAD_REG(I),
										CLK   => CLK,
										RST   => RST,
										DATA  => DATA_IN,
										Q_OUT => BUF_OF_BUFFERS(I,31 DOWNTO 0) -- <= PROBLEM HERE.
									 );
			END GENERATE CASE1;
			
		END GENERATE;
		
END STRUCTURAL; 
										