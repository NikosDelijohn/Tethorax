-- Custom 32 to 1 Generic input Multiplexer.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX32X1 IS

	GENERIC ( INSIZE : INTEGER := 10 );
	
	PORT (
	
			D0 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D1 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D2 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D3 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D4 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D5 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D6 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D7 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D8 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D9 : IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D10: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D11: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D12: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D13: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D14: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D15: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D16: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D17: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D18: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D19: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D20: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D21: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D22: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D23: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D24: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D25: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D26: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D27: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0);
			D28: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D29: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D30: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			D31: IN  STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0) := NULL;
			
			SEL: IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
			
			O  : OUT STD_LOGIC_VECTOR(INSIZE-1 DOWNTO 0)
		);
		
END MUX32X1;

ARCHITECTURE RTL OF MUX32X1 IS

BEGIN

	PROCESS(SEL)
	BEGIN
	
		CASE SEL IS
		    --    OPCODE
			WHEN "00000" => O <= D0;  -- LOADS
			WHEN "00100" => O <= D4;  -- I-OPS
			WHEN "00101" => O <= D5;  -- AUIPC
			WHEN "01000" => O <= D8;  -- STORES
			WHEN "01100" => O <= D12; -- R-OPS
			WHEN "01101" => O <= D13; -- LUI
			WHEN "11000" => O <= D24; -- BRANCHES
			WHEN "11001" => O <= D25; -- JALR
			WHEN "11011" => O <= D27; -- JAL
			WHEN OTHERS  => O <= (OTHERS => 'Z');
		
		END CASE;
		
	END PROCESS;
	
END RTL;
